module pbdebounce(
	input wire clk_1ms,
	input wire button, 
	output reg pbreg
	);
 
	reg [7:0] pbshift;

	always@(posedge clk_1ms) begin
		pbshift=pbshift<<1;// moving to left 2 wei // multiple 2
		pbshift[0]=button;
		if (pbshift==8'b0)
			pbreg=0;
		if (pbshift==8'hFF)// 11111111
			pbreg=1;	
	end
endmodule
// clk_1ms goes through 8 periods,ouput the input
// like pitting off outputing
